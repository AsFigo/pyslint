class gen_c;
  rand bit b;
  
  function pre_randomize();
  endfunction 
  
  function post_randomize();
  endfunction
endclass : gen_c
