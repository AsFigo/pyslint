//----------------------------------------------------
// SPDX-FileCopyrightText: Jayaraman R P,
//                         Verifworks Pvt Ltd,India
// SPDX-License-Identifier: MIT
//----------------------------------------------------
class add;
  bit var1;
  bit var2;

endclass :add 
