//----------------------------------------------------
// SPDX-FileCopyrightText: Srinivasan Venkataramanan,
//                         AsFigo Technologies, UK
// SPDX-License-Identifier: MIT
//----------------------------------------------------

interface af_sv_if ();
  wire  wire_a;
  logic logic_a;
endinterface : af_sv_if

