package pack1;
  import "DPI-C" function int good_dpi_f(input int v, output int o);
  import "DPI-C" function int bad_dpi_f_4st(input integer v, output logic o);
  import "DPI-C" function int bad_dpi_f_4st_1(input integer v, output bit o);
  import "DPI-C" function int bad_dpi_f_4st_def(input v, output o);
endpackage
