//----------------------------------------------------
//----------------------------------------------------
// SPDX-FileCopyrightText: Srinivasan Venkataramanan, 
//                         AsFigo Technologies, UK
// SPDX-License-Identifier: MIT
//----------------------------------------------------

class test_sv_name_chk_30_p_c;
  
endclass : test_sv_name_chk_30_p_c