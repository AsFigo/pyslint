interface af_sv_if;
  import "DPI" function int c_sum();
  import "DPI-C" function logic c_bad_4_st();
  import "DPI-C" function c_bad_implicit_rt();
endinterface : af_sv_if
