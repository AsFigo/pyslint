class gen_c;
  rand bit b;
  
  function void pre_randomize();
  endfunction : pre_randomize 
  
  function void post_randomize();
  endfunction : post_randomize
endclass : gen_c
