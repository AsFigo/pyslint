class gen_c;
  mailbox gbx;
  mailbox #(int) int_mbx;
endclass : gen_c
