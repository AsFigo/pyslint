class add;
  bit var1;
  bit var2;

endclass :add 
