class abstract_ifc #(int cwidth=1, int awidth, int dwidth);
endclass : abstract_ifc

