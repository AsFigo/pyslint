//----------------------------------------------------
// SPDX-FileCopyrightText: Jayaraman R P,
//                         Verifworks Pvt Ltd,India
// SPDX-License-Identifier: MIT
//----------------------------------------------------
class trailing_whitespace;
  bit line_wo_trailing_space;
  bit line_with_trailing_space; 

endclass: trailing_whitespace
