class trailing_whitespace;
  bit line_wo_trailing_space;
  bit line_with_trailing_space; 

endclass: trailing_whitespace
