module empty_loop_f;
    initial
        begin
           for (int i = 0; i < 100; i++) begin
           // empty loop
        end
        end
endmodule