//----------------------------------------------------
//----------------------------------------------------
// SPDX-FileCopyrightText: Mehul Arvind Prajapati
//                         AsFigo Technologies, UK
// SPDX-License-Identifier: MIT
//----------------------------------------------------

class trans_c;
  
endclass : trans_c

class drv_c;

endclass : drv_c
