import "DPI-C"  function dpi_f (bit [3:0] a);

module top ;

endmodule
